module testbech;

bit [7:0] x;
bit enable;
bit clk;
bit rst_n;

bit [254:0][7:0] message = '{181, 25, 235, 188, 90, 218, 170, 64, 253, 234, 223, 250, 224, 247, 139, 115, 151, 34, 135, 27, 243, 0, 83, 95, 240, 25, 70, 184, 81, 195, 120, 136, 11, 76, 89, 70, 192, 10, 229, 6, 241, 217, 206, 199, 198, 116, 115, 147, 133, 65, 89, 112, 105, 158, 70, 97, 177, 189, 207, 151, 231, 55, 241, 192, 164, 145, 144, 217, 250, 71, 135, 4, 210, 214, 170, 24, 12, 8, 106, 100, 171, 44, 169, 158, 52, 157, 72, 51, 176, 163, 189, 68, 60, 147, 177, 92, 186, 80, 12, 18, 16, 103, 4, 70, 211, 136, 24, 251, 14, 152, 57, 205, 218, 242, 203, 51, 149, 127, 159, 227, 161, 143, 73, 101, 152, 193, 223, 43, 190, 113, 185, 87, 129, 80, 253, 35, 176, 38, 195, 207, 159, 95, 117, 220, 254, 50, 149, 126, 215, 75, 40, 185, 192, 178, 247, 220, 36, 239, 233, 121, 166, 56, 12, 113, 100, 54, 13, 142, 14, 183, 231, 96, 44, 166, 98, 128, 156, 204, 180, 220, 147, 55, 150, 11, 74, 192, 67, 112, 77, 113, 169, 122, 65, 64, 59, 176, 144, 95, 16, 203, 106, 83, 242, 144, 243, 97, 103, 226, 88, 205, 248, 62, 226, 140, 200, 50, 233, 220, 189, 134, 230, 240, 214,
94, 53, 240, 154, 218, 166, 92, 205, 3, 237, 80, 173, 136, 175, 240, 66, 2, 99, 119, 162, 54, 251, 135, 217, 187, 197, 10, 60, 135, 217, 191, 90};




rsdec u_rsdec (
    .x              (x),
    .error          (),
    .with_error     (),
    .enable         (enable),
    .valid          (),
    .k              (32),
    .clk            (clk),
    .rst_n          (rst_n)
);

bit [7:0] a, b;

gf_mul u_gf_mul (
    .a(a),
    .b(b),
    .z()
);


gf_mul_lut u_gf_mul_lut (
    .a(a),
    .b(b),
    .z()
);

initial begin
    a = 30;
    b = 140;
    #20
    a = 52;
    b = 101;
    #20
    a = 240;
    b = 14;
    #20
    a = 18;
    b = 197;
    #20
    a = 0;
    b = 197;
    #20
    a = 18;
    b = 0;
end


initial begin
    clk <= 0;
    forever #10 clk <= ~clk;
end

initial begin
    x <= 0;
    enable <= 0;
    rst_n <= 0;
    repeat(5) @(posedge clk);
    rst_n <= 1;

    repeat(5) @(posedge clk);

    enable <= 1;
    for (int i=254; i >=0; i--) begin
        x <= message[i];
        @(posedge clk);
    end

end

endmodule
